CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 3 100 10
176 80 1364 707
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 0 0
20 Package,Description,
42 C:\Program Files\CircuitMaker 2000\BOM.DAT
0 7
0 4 0.500000 0.500000
344 176 457 273
9437202 0
0
6 Title:
5 Name:
0
0
0
12
13 Logic Switch~
5 83 360 0 10 11
0 17 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 V3
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
4484 0 0
2
5.89884e-315 0
0
7 Ground~
168 721 28 0 1 3
0 2
0
0 0 53360 0
0
4 GND1
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
5996 0 0
2
5.89884e-315 0
0
9 2-In AND~
219 662 251 0 3 22
0 15 11 14
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 U4B
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 3 0
1 U
7804 0 0
2
5.89884e-315 0
0
9 2-In AND~
219 484 242 0 3 22
0 13 12 15
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 U4A
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 3 0
1 U
5523 0 0
2
5.89884e-315 0
0
2 +V
167 837 328 0 1 3
0 18
0
0 0 54256 270
2 5V
-7 -15 7 -7
2 V2
-7 -25 7 -17
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
3330 0 0
2
5.89884e-315 0
0
7 Pulser~
4 89 424 0 10 12
0 19 20 21 16 0 0 5 5 5
7
0
0 0 4656 0
0
2 V1
-7 -28 7 -20
0
0
0
0
0
4 SIP2
9

0 1 2 3 4 1 2 3 4 0
0 0 0 512 1 0 0 0
1 V
3465 0 0
2
5.89884e-315 0
0
6 74112~
219 718 355 0 7 32
0 18 14 16 14 18 22 10
0
0 0 4720 0
5 74112
4 -60 39 -52
3 U3B
22 -61 43 -53
0
15 DVCC=16;DGND=8;
73 %D [%16bi %8bi %1i %2i %3i %4i %5i][%16bo %1o %2o %3o %4o %5o %6o %7o] %M
0
12 type:digital
5 DIP16
32

0 10 11 13 12 14 7 9 4 3
1 2 15 6 5 10 11 13 12 14
7 9 0 0 0 0 0 0 0 0
0 0 0
65 0 0 512 2 2 2 0
1 U
8396 0 0
2
5.89884e-315 0
0
6 74112~
219 571 355 0 7 32
0 18 15 16 15 18 23 11
0
0 0 4720 0
5 74112
4 -60 39 -52
3 U3A
22 -61 43 -53
0
15 DVCC=16;DGND=8;
73 %D [%16bi %8bi %1i %2i %3i %4i %5i][%16bo %1o %2o %3o %4o %5o %6o %7o] %M
0
12 type:digital
5 DIP16
32

0 4 3 1 2 15 6 5 4 3
1 2 15 6 5 10 11 13 12 14
7 9 0 0 0 0 0 0 0 0
0 0 0
65 0 0 512 2 1 2 0
1 U
3685 0 0
2
5.89883e-315 0
0
6 74112~
219 412 355 0 7 32
0 18 13 16 13 18 24 12
0
0 0 4720 0
5 74112
4 -60 39 -52
3 U2B
22 -61 43 -53
0
15 DVCC=16;DGND=8;
73 %D [%16bi %8bi %1i %2i %3i %4i %5i][%16bo %1o %2o %3o %4o %5o %6o %7o] %M
0
12 type:digital
5 DIP16
32

0 10 11 13 12 14 7 9 4 3
1 2 15 6 5 10 11 13 12 14
7 9 0 0 0 0 0 0 0 0
0 0 0
65 0 0 512 2 2 1 0
1 U
7849 0 0
2
5.89883e-315 0
0
6 74112~
219 261 355 0 7 32
0 18 17 16 17 18 25 13
0
0 0 4720 0
5 74112
4 -60 39 -52
3 U2A
22 -61 43 -53
0
15 DVCC=16;DGND=8;
73 %D [%16bi %8bi %1i %2i %3i %4i %5i][%16bo %1o %2o %3o %4o %5o %6o %7o] %M
0
12 type:digital
5 DIP16
32

0 4 3 1 2 15 6 5 4 3
1 2 15 6 5 10 11 13 12 14
7 9 0 0 0 0 0 0 0 0
0 0 0
65 0 0 512 2 1 1 0
1 U
6343 0 0
2
5.89883e-315 0
0
6 74LS48
188 405 135 0 14 29
0 10 11 12 13 26 27 9 8 7
6 5 4 3 28
0
0 0 4848 0
7 74LS248
-24 -60 25 -52
2 U1
-7 -61 7 -53
0
15 DVCC=16;DGND=8;
119 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %14i]
+ [%16bo %1o %2o %3o %4o %5o %6o %14o %7o %8o %9o %10o %11o %12o %13o] %M
0
12 type:digital
5 DIP16
29

0 6 2 1 7 3 5 14 15 9
10 11 12 13 4 6 2 1 7 3
5 14 15 9 10 11 12 13 4 0
65 0 0 512 1 0 0 0
1 U
7376 0 0
2
5.89883e-315 0
0
9 CC 7-Seg~
183 742 78 0 17 19
10 3 4 5 6 7 8 9 29 2
0 0 0 1 1 0 1 2
0
0 0 21104 0
7 AMBERCC
9 -41 58 -33
5 DISP1
30 -4 65 4
0
0
32 %D %1 %2 %3 %4 %5 %6 %7 %8 %9 %S
0
0
0
19

0 1 2 3 4 5 6 7 8 9
1 2 3 4 5 6 7 8 9 0
88 0 0 512 1 0 0 0
4 DISP
9156 0 0
2
5.89883e-315 0
0
36
1 9 2 0 0 4224 0 2 12 0 0 3
721 22
742 22
742 36
13 1 3 0 0 12416 0 11 12 0 0 5
437 153
528 153
528 194
721 194
721 114
12 2 4 0 0 12416 0 11 12 0 0 5
437 144
540 144
540 184
727 184
727 114
11 3 5 0 0 12416 0 11 12 0 0 5
437 135
551 135
551 173
733 173
733 114
10 4 6 0 0 12416 0 11 12 0 0 5
437 126
564 126
564 158
739 158
739 114
9 5 7 0 0 12416 0 11 12 0 0 5
437 117
576 117
576 147
745 147
745 114
8 6 8 0 0 12416 0 11 12 0 0 5
437 108
589 108
589 136
751 136
751 114
7 7 9 0 0 4224 0 11 12 0 0 5
437 99
599 99
599 123
757 123
757 114
7 1 10 0 0 8320 0 7 11 0 0 5
742 319
742 204
367 204
367 99
373 99
7 2 11 0 0 8320 0 8 11 0 0 5
595 319
595 222
333 222
333 108
373 108
7 3 12 0 0 8320 0 9 11 0 0 5
436 319
436 238
308 238
308 117
373 117
7 4 13 0 0 4224 0 10 11 0 0 3
285 319
285 126
373 126
4 3 14 0 0 8320 0 7 3 0 0 3
694 337
683 337
683 251
3 2 14 0 0 0 0 3 7 0 0 3
683 251
683 319
694 319
2 7 11 0 0 0 0 3 8 0 0 4
638 260
622 260
622 319
595 319
1 3 15 0 0 4224 0 3 4 0 0 2
638 242
505 242
4 0 15 0 0 0 0 8 0 0 18 3
547 337
521 337
521 319
3 2 15 0 0 0 0 4 8 0 0 3
505 242
505 319
547 319
4 0 13 0 0 0 0 9 0 0 20 3
388 337
357 337
357 318
0 7 13 0 0 0 0 0 10 21 0 3
357 318
357 319
285 319
1 2 13 0 0 0 0 4 9 0 0 4
460 233
357 233
357 319
388 319
2 7 12 0 0 0 0 4 9 0 0 3
460 251
460 319
436 319
3 0 16 0 0 4096 0 10 0 0 26 2
231 328
231 395
3 0 16 0 0 0 0 9 0 0 26 2
382 328
382 395
3 0 16 0 0 0 0 8 0 0 26 2
541 328
541 395
4 3 16 0 0 12416 0 6 7 0 0 5
119 424
231 424
231 395
688 395
688 328
1 0 17 0 0 4224 0 1 0 0 28 4
95 360
185 360
185 327
200 327
4 2 17 0 0 0 0 10 10 0 0 4
237 337
200 337
200 319
237 319
5 5 18 0 0 4096 0 9 10 0 0 2
412 367
261 367
5 5 18 0 0 4224 0 8 9 0 0 2
571 367
412 367
5 5 18 0 0 0 0 7 8 0 0 2
718 367
571 367
1 5 18 0 0 0 0 5 7 0 0 3
825 327
825 367
718 367
1 1 18 0 0 0 0 7 5 0 0 3
718 292
825 292
825 327
1 1 18 0 0 0 0 8 7 0 0 2
571 292
718 292
1 1 18 0 0 0 0 9 8 0 0 2
412 292
571 292
1 1 18 0 0 0 0 10 9 0 0 2
261 292
412 292
1
-24 0 0 0 400 0 0 0 0 3 2 1 34
14 Century Gothic
0 0 0 25
14 25 400 65
24 33 389 63
25 4-BIT SYNCHRONOUS COUNTER
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
